module LED(
	input sw,
	output LED

);

assign LED = sw;

endmodule
